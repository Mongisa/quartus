module lut1(A,Y);
input wire [4:0] A;
output reg Y;

//Mintermini
/*assign Y = 
	(~(A[4] | A[3] | A[2] | A[1]) & A[0]) | //m1
	(~(A[4] | A[3] | A[2] | A[0]) & A[1]) | //m2
	(~(A[4] | A[3] | A[2]) & A[1] & A[0]) | //m3
	(~(A[4] | A[3] | A[1] | A[0]) & A[2]) | //m4
	(~(A[4] | A[3] | A[0]) & A[2] & A[1]) | //m6
	(~(A[4] | A[2] | A[1] | A[0]) & A[3]) | //m8
	(~(A[4] | A[2] | A[0]) & A[3] & A[1]) | //m10
	(~(A[4] | A[2]) & A[3] & A[1] & A[0]) | //m11
	(~(A[4] | A[0]) & A[3] & A[2] & A[1]) | //m14
	(~(A[3] | A[2] | A[1]) & A[4] & A[0]) | //m17
	(~(A[3] | A[2] | A[0]) & A[4] & A[1]) | //m18
	(~(A[3] | A[1]) & A[4] & A[2] & A[0]) | //m21
	(A[4] & ~A[3] & A[2] & A[1] & ~A[0]) | //m22
	(A[4] & ~A[3] & A[2] & A[1] & A[0]) | //m23
	(A[4] & A[3] & ~A[2] & ~A[1] & ~A[0]) | //m24
	(A[4] & A[3] & ~A[2] & ~A[1] & A[0]) | //m25
	(A[4] & A[3] & ~A[2] & A[1] & A[0]) | //m27
	(A[4] & A[3] & A[2] & ~A[1] & ~A[0]) | //m28
	(A[4] & A[3] & A[2] & ~A[1] & A[0]) | //m29
	(A[4] & A[3] & A[2] & A[1] & ~A[0]); //m30*/

//Blocco procedurale
always @ (A)
begin
	case (A)
		5'd0: Y<=1'b0;
		5'd5: Y<=1'b0;
		5'd7: Y<=1'b0;
		5'd9: Y<=1'b0;
		5'd12: Y<=1'b0;
		5'd13: Y<=1'b0;
		5'd15: Y<=1'b0;
		5'd16: Y<=1'b0;
		5'd19: Y<=1'b0;
		5'd20: Y<=1'b0;
		5'd26: Y<=1'b0;
		5'd31: Y<=1'b0;
		default: Y<=1'b1;
	endcase
end
endmodule