module seven_seg_decoder(A,Y);
input wire [3:0] A;
output reg [6:0] Y;

always@(A)
begin
	case (A)
	4'd0: Y<= 7'b100_0000; //0
	4'd1: Y<= 7'b111_1001; //1
	4'd2: Y<= 7'b010_0100; //2
	4'd3: Y<= 7'b011_0000; //3
	4'd4: Y<= 7'b001_1001; //4
	4'd5: Y<= 7'b001_0010; //5
	4'd6: Y<= 7'b000_0010; //6
	4'd7: Y<= 7'b101_1000; //7
	4'd8: Y<= 7'b000_0000; //8
	4'd9: Y<= 7'b001_0000; //9
	4'd10: Y<= 7'b000_1000; //10 (A)
	4'd11: Y<= 7'b000_0011; //11 (B)
	4'd12: Y<= 7'b100_0110; //12 (C)
	4'd13: Y<= 7'b010_0001; //13 (D)
	4'd14: Y<= 7'b000_0110; //14 (E)
	4'd15: Y<= 7'b000_1110; //15 (F)
	default: Y<= 7'd0;
	endcase
end
endmodule